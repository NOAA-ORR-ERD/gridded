netcdf fvcom.nc {
dimensions:
        nele = 36477 ;
        node = 20689 ;
        siglay = 6 ;
        siglev = 7 ;
        three = 3 ;
        time = UNLIMITED ; // (24 currently)
        DateStrLen = 26 ;
variables:
        int nprocs ;
                nprocs:long_name = "number of processors" ;
        int partition(nele) ;
                partition:long_name = "partition" ;
        float x(node) ;
                x:long_name = "nodal x-coordinate" ;
                x:units = "meters" ;
        float y(node) ;
                y:long_name = "nodal y-coordinate" ;
                y:units = "meters" ;
        float lon(node) ;
                lon:long_name = "nodal longitude" ;
                lon:standard_name = "longitude" ;
                lon:units = "degrees_east" ;
        float lat(node) ;
                lat:long_name = "nodal latitude" ;
                lat:standard_name = "latitude" ;
                lat:units = "degrees_north" ;
        float xc(nele) ;
                xc:long_name = "zonal x-coordinate" ;
                xc:units = "meters" ;
        float yc(nele) ;
                yc:long_name = "zonal y-coordinate" ;
                yc:units = "meters" ;
        float lonc(nele) ;
                lonc:long_name = "zonal longitude" ;
                lonc:standard_name = "longitude" ;
                lonc:units = "degrees_east" ;
        float latc(nele) ;
                latc:long_name = "zonal latitude" ;
                latc:standard_name = "latitude" ;
                latc:units = "degrees_north" ;
        float siglay(siglay, node) ;
                siglay:long_name = "Sigma Layers" ;
                siglay:standard_name = "ocean_sigma/general_coordinate" ;
                siglay:positive = "up" ;
                siglay:valid_min = -1.f ;
                siglay:valid_max = 0.f ;
                siglay:formula_terms = "sigma: siglay eta: zeta depth: h" ;
        float siglev(siglev, node) ;
                siglev:long_name = "Sigma Levels" ;
                siglev:standard_name = "ocean_sigma/general_coordinate" ;
                siglev:positive = "up" ;
                siglev:valid_min = -1.f ;
                siglev:valid_max = 0.f ;
                siglev:formula_terms = "sigma:siglay eta: zeta depth: h" ;
        float siglay_center(siglay, nele) ;
                siglay_center:long_name = "Sigma Layers" ;
                siglay_center:standard_name = "ocean_sigma/general_coordinate" ;
                siglay_center:positive = "up" ;
                siglay_center:valid_min = -1.f ;
                siglay_center:valid_max = 0.f ;
                siglay_center:formula_terms = "sigma: siglay_center eta: zeta_center depth: h_center" ;
        float siglev_center(siglev, nele) ;
                siglev_center:long_name = "Sigma Levels" ;
                siglev_center:standard_name = "ocean_sigma/general_coordinate" ;
                siglev_center:positive = "up" ;
                siglev_center:valid_min = -1.f ;
                siglev_center:valid_max = 0.f ;
                siglev_center:formula_terms = "sigma:siglay_center eta: zeta_center depth: h_center" ;
        float h_center(nele) ;
                h_center:long_name = "Bathymetry" ;
                h_center:standard_name = "sea_floor_depth_below_geoid" ;
                h_center:units = "m" ;
                h_center:positive = "down" ;
                h_center:grid = "grid1 grid3" ;
                h_center:coordinates = "latc lonc" ;
                h_center:grid_location = "center" ;
        float h(node) ;
                h:long_name = "Bathymetry" ;
                h:standard_name = "sea_floor_depth_below_geoid" ;
                h:units = "m" ;
                h:positive = "down" ;
                h:grid = "Bathymetry_Mesh" ;
                h:coordinates = "lat lon" ;
                h:type = "data" ;
        int nv(three, nele) ;
                nv:long_name = "nodes surrounding element" ;
        int iint(time) ;
                iint:long_name = "internal mode iteration number" ;
        float time(time) ;
                time:long_name = "time" ;
                time:units = "days since 1970-01-01 00:00:00" ;
                time:format = "defined reference date" ;
                time:time_zone = "UTC" ;
        int Itime(time) ;
                Itime:units = "days since 1970-01-01 00:00:00" ;
                Itime:format = "defined reference date" ;
                Itime:time_zone = "UTC" ;
        int Itime2(time) ;
                Itime2:units = "msec since 00:00:00" ;
                Itime2:time_zone = "UTC" ;
        char Times(time, DateStrLen) ;
                Times:time_zone = "UTC" ;
        float zeta(time, node) ;
                zeta:long_name = "Water Surface Elevation" ;
                zeta:units = "meters" ;
                zeta:positive = "up" ;
                zeta:standard_name = "sea_surface_height_above_geoid" ;
                zeta:grid = "Bathymetry_Mesh" ;
                zeta:coordinates = "time lat lon" ;
                zeta:type = "data" ;
                zeta:location = "node" ;
        float u(time, siglay, nele) ;
                u:long_name = "Eastward Water Velocity" ;
                u:standard_name = "eastward_sea_water_velocity" ;
                u:units = "meters s-1" ;
                u:grid = "fvcom_grid" ;
                u:type = "data" ;
                u:coordinates = "time siglay latc lonc" ;
                u:mesh = "fvcom_mesh" ;
                u:location = "face" ;
        float v(time, siglay, nele) ;
                v:long_name = "Northward Water Velocity" ;
                v:standard_name = "Northward_sea_water_velocity" ;
                v:units = "meters s-1" ;
                v:grid = "fvcom_grid" ;
                v:type = "data" ;
                v:coordinates = "time siglay latc lonc" ;
                v:mesh = "fvcom_mesh" ;
                v:location = "face" ;
        float tauc(time, nele) ;
                tauc:long_name = "bed stress magnitude from currents" ;
                tauc:note1 = "this stress is bottom boundary condtion on velocity field" ;
                tauc:note2 = "dimensions are stress/rho" ;
                tauc:units = "m^2 s^-2" ;
                tauc:grid = "fvcom_grid" ;
                tauc:type = "data" ;
                tauc:coordinates = "time latc lonc" ;
                tauc:mesh = "fvcom_mesh" ;
                tauc:location = "face" ;
        float temp(time, siglay, node) ;
                temp:long_name = "temperature" ;
                temp:standard_name = "sea_water_temperature" ;
                temp:units = "degrees_C" ;
                temp:grid = "fvcom_grid" ;
                temp:coordinates = "time siglay lat lon" ;
                temp:type = "data" ;
                temp:mesh = "fvcom_mesh" ;
                temp:location = "node" ;
        float salinity(time, siglay, node) ;
                salinity:long_name = "salinity" ;
                salinity:standard_name = "sea_water_salinity" ;
                salinity:units = "1e-3" ;
                salinity:grid = "fvcom_grid" ;
                salinity:coordinates = "time siglay lat lon" ;
                salinity:type = "data" ;
                salinity:mesh = "fvcom_mesh" ;
                salinity:location = "node" ;
        float short_wave(time, node) ;
                short_wave:long_name = "Short Wave Radiation" ;
                short_wave:units = "W m-2" ;
                short_wave:grid = "fvcom_grid" ;
                short_wave:coordinates = "time lat lon" ;
                short_wave:type = "data" ;
                short_wave:mesh = "fvcom_mesh" ;
                short_wave:location = "node" ;
        float net_heat_flux(time, node) ;
                net_heat_flux:long_name = "Surface Net Heat Flux" ;
                net_heat_flux:units = "W m-2" ;
                net_heat_flux:grid = "fvcom_grid" ;
                net_heat_flux:coordinates = "time lat lon" ;
                net_heat_flux:type = "data" ;
                net_heat_flux:mesh = "fvcom_mesh" ;
                net_heat_flux:location = "node" ;
        float sensible_heat_flux(time, node) ;
                sensible_heat_flux:long_name = "Sensible Heat Flux" ;
                sensible_heat_flux:units = "W m-2" ;
                sensible_heat_flux:grid = "fvcom_grid" ;
                sensible_heat_flux:coordinates = "time lat lon" ;
                sensible_heat_flux:type = "data" ;
                sensible_heat_flux:mesh = "fvcom_mesh" ;
                sensible_heat_flux:location = "node" ;
        float latent_heat_flux(time, node) ;
                latent_heat_flux:long_name = "Latent Heat Flux" ;
                latent_heat_flux:units = "W m-2" ;
                latent_heat_flux:grid = "fvcom_grid" ;
                latent_heat_flux:coordinates = "time lat lon" ;
                latent_heat_flux:type = "data" ;
                latent_heat_flux:mesh = "fvcom_mesh" ;
                latent_heat_flux:location = "node" ;
        float long_wave(time, node) ;
                long_wave:long_name = "Long Wave Radiation" ;
                long_wave:units = "W m-2" ;
                long_wave:grid = "fvcom_grid" ;
                long_wave:coordinates = "time lat lon" ;
                long_wave:type = "data" ;
                long_wave:mesh = "fvcom_mesh" ;
                long_wave:location = "node" ;
        float uwind_speed(time, nele) ;
                uwind_speed:long_name = "Eastward Wind Velocity" ;
                uwind_speed:standard_name = "eastward wind" ;
                uwind_speed:units = "meters s-1" ;
                uwind_speed:grid = "fvcom_grid" ;
                uwind_speed:coordinates = "time latc lonc" ;
                uwind_speed:type = "data" ;
                uwind_speed:mesh = "fvcom_mesh" ;
                uwind_speed:location = "face" ;
        float vwind_speed(time, nele) ;
                vwind_speed:long_name = "Northward Wind Velocity" ;
                vwind_speed:standard_name = "northward wind" ;
                vwind_speed:units = "meters s-1" ;
                vwind_speed:grid = "fvcom_grid" ;
                vwind_speed:coordinates = "time latc lonc" ;
                vwind_speed:type = "data" ;
                vwind_speed:mesh = "fvcom_mesh" ;
                vwind_speed:location = "face" ;
        int wet_nodes(time, node) ;
                wet_nodes:long_name = "Wet_Nodes" ;
                wet_nodes:grid = "fvcom_grid" ;
                wet_nodes:type = "data" ;
                wet_nodes:coordinates = "time lat lon" ;
                wet_nodes:mesh = "fvcom_mesh" ;
                wet_nodes:location = "node" ;
        int wet_cells(time, nele) ;
                wet_cells:long_name = "Wet_Cells" ;
                wet_cells:grid = "fvcom_grid" ;
                wet_cells:type = "data" ;
                wet_cells:coordinates = "time latc lonc" ;
                wet_cells:mesh = "fvcom_mesh" ;
                wet_cells:location = "face" ;
        int wet_nodes_prev_int(time, node) ;
                wet_nodes_prev_int:long_name = "Wet_Nodes_At_Previous_Internal_Step" ;
                wet_nodes_prev_int:grid = "fvcom_grid" ;
                wet_nodes_prev_int:type = "data" ;
                wet_nodes_prev_int:coordinates = "time lat lon" ;
                wet_nodes_prev_int:mesh = "fvcom_mesh" ;
                wet_nodes_prev_int:location = "node" ;
        int wet_cells_prev_int(time, nele) ;
                wet_cells_prev_int:long_name = "Wet_Cells_At_Previous_Internal_Step" ;
                wet_cells_prev_int:grid = "fvcom_grid" ;
                wet_cells_prev_int:type = "data" ;
                wet_cells_prev_int:coordinates = "time latc lonc" ;
                wet_cells_prev_int:mesh = "fvcom_mesh" ;
                wet_cells_prev_int:location = "face" ;
        int wet_cells_prev_ext(time, nele) ;
                wet_cells_prev_ext:long_name = "Wet_Cells_At_Previous_External_Step" ;
                wet_cells_prev_ext:grid = "fvcom_grid" ;
                wet_cells_prev_ext:type = "data" ;
        float aice(time, node) ;
                aice:long_name = "ice area" ;
                aice:standard_name = "ice_area_category" ;
                aice:units = "" ;
                aice:grid = "fvcom_grid" ;
                aice:coordinates = "lat lon" ;
                aice:type = "data" ;
        float vice(time, node) ;
                vice:long_name = "ice volume per unit grid area" ;
                vice:standard_name = "ice_volume_category" ;
                vice:units = "m" ;
                vice:grid = "fvcom_grid" ;
                vice:coordinates = "lat lon" ;
                vice:type = "data" ;
        float tsfc(time, node) ;
                tsfc:long_name = "ice surface temperature" ;
                tsfc:standard_name = "ice_surface_temperature" ;
                tsfc:units = "deg C" ;
                tsfc:grid = "fvcom_grid" ;
                tsfc:coordinates = "lat lon" ;
                tsfc:type = "data" ;
        float uuice(time, nele) ;
                uuice:long_name = "Ice x-velocity" ;
                uuice:units = "meters s-1" ;
                uuice:grid = "fvcom_grid" ;
                uuice:type = "data" ;
        float vvice(time, nele) ;
                vvice:long_name = "Ice y-velocity" ;
                vvice:units = "meters s-1" ;
                vvice:grid = "fvcom_grid" ;
                vvice:type = "data" ;

// global attributes:
                :title = "Huron Erie Connecting Waterways version \"\". Forecast Run \"031400\". 2023-03-14 00" ;
                :institution = "School for Marine Science and Technology" ;
                :source = "FVCOM_4.3" ;
                :history = "model started at: 14/03/2023   05:41" ;
                :references = "http://fvcom.smast.umassd.edu, http://codfish.smast.umassd.edu" ;
                :Conventions = "CF-1.0" ;
                :CoordinateSystem = "GeoReferenced" ;
                :CoordinateProjection = "lonlat" ;
                :Tidal_Forcing = "Tidal Forcing Time Series Title: UNKNOWN" ;
                :River_Forcing = "THERE ARE 8 RIVERS IN THIS MODEL.\n",
                        "RIVER INFLOW IS ON THE nodes WHERE TEMPERATURE AND SALINITY ARE specified IN THE MODEL.\n",
                        "THE FOLLOWING RIVER NAMES ARE USED:\n",
                        "BlackRiver01\n",
                        "PineRiver01\n",
                        "BelleRiver01\n",
                        "SydenhamRiver01\n",
                        "ClintonRiver01\n",
                        "ClintonCutoff01\n",
                        "ThamesRiver01\n",
                        "RiverRouge01" ;
                :GroundWater_Forcing = "GROUND WATER FORCING IS OFF!" ;
                :Surface_Heat_Forcing = "FVCOM variable surface heat forcing file:\n",
                        "FILE NAME:031400_met.nc\n",
                        "SOURCE:FVCOM grid (unstructured) surface forcing\n",
                        "Unknown start date meta data format" ;
                :Surface_Wind_Forcing = "FVCOM variable surface Wind forcing:\n",
                        "FILE NAME:031400_met.nc\n",
                        "SOURCE:FVCOM grid (unstructured) surface forcing\n",
                        "Unknown start date meta data format" ;
                :Surface_PrecipEvap_Forcing = "SURFACE PRECIPITATION FORCING IS OFF" ;
                :Ice_Model_Forcing = "FVCOM variable surface ice model forcing:\n",
                        "FILE NAME:031400_met.nc\n",
                        "SOURCE:FVCOM grid (unstructured) surface forcing\n",
                        "Unknown start date meta data format" ;
}