netcdf TBOFS_wind_test {
dimensions:
        time = UNLIMITED ; // (49 currently)
        eta_rho = 145 ;
        xi_rho = 176 ;
        eta_psi = 144 ;
        xi_psi = 175 ;
        eta_u = 145 ;
        xi_u = 175 ;
        eta_v = 144 ;
        xi_v = 176 ;
variables:
        float time(time) ;
                time:units = "hours since 2023-03-12 18:00:00.000 UTC" ;
        double lon_rho(eta_rho, xi_rho) ;
                lon_rho:units = "degrees_east" ;
                lon_rho:long_name = "longitude of RHO-points" ;
                lon_rho:standard_name = "longitude" ;
                lon_rho:field = "longitude" ;
                lon_rho:_CoordinateAxisType = "Lon" ;
        double lat_rho(eta_rho, xi_rho) ;
                lat_rho:units = "degrees_north" ;
                lat_rho:long_name = "latitude of RHO-points" ;
                lat_rho:standard_name = "latitude" ;
                lat_rho:field = "latitude" ;
                lat_rho:_CoordinateAxisType = "Lat" ;
        double mask_rho(eta_rho, xi_rho) ;
                mask_rho:long_name = "mask on RHO-points" ;
                mask_rho:standard_name = "land_sea_mask_at_cell_center" ;
                mask_rho:flag_values = 0., 1. ;
                mask_rho:flag_meanings = "land water" ;
                mask_rho:grid = "grid" ;
                mask_rho:location = "face" ;
                mask_rho:coordinates = "lat_rho lon_rho " ;
        double lon_psi(eta_psi, xi_psi) ;
                lon_psi:units = "degrees_east" ;
                lon_psi:long_name = "longitude of PSI-points" ;
                lon_psi:standard_name = "longitude" ;
                lon_psi:field = "longitude" ;
                lon_psi:_CoordinateAxisType = "Lon" ;
        double lat_psi(eta_psi, xi_psi) ;
                lat_psi:units = "degrees_north" ;
                lat_psi:long_name = "latitude of PSI-points" ;
                lat_psi:standard_name = "latitude" ;
                lat_psi:field = "latitude" ;
                lat_psi:_CoordinateAxisType = "Lat" ;
        double mask_psi(eta_psi, xi_psi) ;
                mask_psi:long_name = "mask on psi-points" ;
                mask_psi:standard_name = "land_sea_mask_at_cell_corners" ;
                mask_psi:flag_values = 0., 1. ;
                mask_psi:flag_meanings = "land water" ;
                mask_psi:grid = "grid" ;
                mask_psi:location = "node" ;
                mask_psi:coordinates = "lat_psi lon_psi " ;
        double lon_u(eta_u, xi_u) ;
                lon_u:units = "degrees_east" ;
                lon_u:long_name = "longitude of U-points" ;
                lon_u:standard_name = "longitude" ;
                lon_u:field = "longitude" ;
                lon_u:_CoordinateAxisType = "Lon" ;
        double lat_u(eta_u, xi_u) ;
                lat_u:units = "degrees_north" ;
                lat_u:long_name = "latitude of U-points" ;
                lat_u:standard_name = "latitude" ;
                lat_u:field = "latitude" ;
                lat_u:_CoordinateAxisType = "Lat" ;
        double mask_u(eta_u, xi_u) ;
                mask_u:long_name = "mask on U-points" ;
                mask_u:standard_name = "land_sea_mask_at_cell_y_edges" ;
                mask_u:flag_values = 0., 1. ;
                mask_u:flag_meanings = "land water" ;
                mask_u:grid = "grid" ;
                mask_u:location = "edge1" ;
                mask_u:coordinates = "lat_u lon_u " ;
        double lon_v(eta_v, xi_v) ;
                lon_v:units = "degrees_east" ;
                lon_v:long_name = "longitude of V-points" ;
                lon_v:standard_name = "longitude" ;
                lon_v:field = "longitude" ;
                lon_v:_CoordinateAxisType = "Lon" ;
        double lat_v(eta_v, xi_v) ;
                lat_v:units = "degrees_north" ;
                lat_v:long_name = "latitude of V-points" ;
                lat_v:standard_name = "latitude" ;
                lat_v:field = "latitude" ;
                lat_v:_CoordinateAxisType = "Lat" ;
        float Uwind(time, eta_rho, xi_rho) ;
                Uwind:units = "meter second-1" ;
                Uwind:long_name = "surface u-wind component" ;
                Uwind:standard_name = "grid_eastward_wind" ;
                Uwind:time = "ocean_time" ;
                Uwind:cell_methods = "ocean_time: point" ;
                Uwind:grid = "grid" ;
                Uwind:location = "face" ;
                Uwind:coordinates = "time_run time lat_rho lon_rho " ;
                Uwind:field = "u-wind" ;
        float Vwind(time, eta_rho, xi_rho) ;
                Vwind:units = "meter second-1" ;
                Vwind:long_name = "surface v-wind component" ;
                Vwind:standard_name = "grid_northward_wind" ;
                Vwind:time = "ocean_time" ;
                Vwind:cell_methods = "ocean_time: point" ;
                Vwind:grid = "grid" ;
                Vwind:location = "face" ;
                Vwind:coordinates = "time_run time lat_rho lon_rho " ;
                Vwind:field = "v-wind" ;
}