netcdf wcofs_fc {
dimensions:
	ocean_time = UNLIMITED ; // (24 currently)
	eta_rho = 205 ;
	xi_rho = 348 ;
	eta_psi = 204 ;
	xi_psi = 347 ;
	eta_u = 205 ;
	xi_u = 347 ;
	eta_v = 204 ;
	xi_v = 348 ;
variables:
	float ocean_time(ocean_time) ;
		ocean_time:units = "seconds since 2016-01-01 00:00:00" ;
		ocean_time:cell_methods = "ocean_time: mean" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
		lon_rho:field = "lon_rho, scalar" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
		lat_rho:field = "lat_rho, scalar" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:flag_values = 0., 1. ;
		mask_rho:flag_meanings = "land water" ;
		mask_rho:grid = "grid" ;
		mask_rho:location = "face" ;
		mask_rho:coordinates = "lon_rho lat_rho" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
		lon_psi:standard_name = "longitude" ;
		lon_psi:field = "lon_psi, scalar" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
		lat_psi:standard_name = "latitude" ;
		lat_psi:field = "lat_psi, scalar" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on psi-points" ;
		mask_psi:flag_values = 0., 1. ;
		mask_psi:flag_meanings = "land water" ;
		mask_psi:grid = "grid" ;
		mask_psi:location = "node" ;
		mask_psi:coordinates = "lon_psi lat_psi" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:standard_name = "longitude" ;
		lon_u:field = "lon_u, scalar" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:standard_name = "latitude" ;
		lat_u:field = "lat_u, scalar" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:flag_values = 0., 1. ;
		mask_u:flag_meanings = "land water" ;
		mask_u:grid = "grid" ;
		mask_u:location = "edge1" ;
		mask_u:coordinates = "lon_u lat_u" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:standard_name = "longitude" ;
		lon_v:field = "lon_v, scalar" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:standard_name = "latitude" ;
		lat_v:field = "lat_v, scalar" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:flag_values = 0., 1. ;
		mask_v:flag_meanings = "land water" ;
		mask_v:grid = "grid" ;
		mask_v:location = "edge2" ;
		mask_v:coordinates = "lon_v lat_v" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between XI-axis and EAST" ;
		angle:units = "radians" ;
		angle:grid = "grid" ;
		angle:location = "face" ;
		angle:coordinates = "lon_rho lat_rho" ;
		angle:field = "angle, scalar" ;
	float u(ocean_time, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:grid = "grid" ;
		u:location = "edge1" ;
		u:coordinates = "lon_u lat_u " ;
		u:field = "u-velocity, scalar, series" ;
		u:cell_methods = "ocean_time: mean" ;
	float v(ocean_time, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:grid = "grid" ;
		v:location = "edge2" ;
		v:coordinates = "lon_v lat_v " ;
		v:field = "v-velocity, scalar, series" ;
		v:cell_methods = "ocean_time: mean" ;

// global attributes:
		:history = "Wed Apr  6 14:39:04 2022: ncra -Y ncrcat wcofs_fc.nc" ;
		:NCO = "netCDF Operators version 5.0.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:nco_input_file_number = 24 ;
		:nco_input_file_list = "wcofs_20220406_t03z_f003.nc wcofs_20220406_t03z_f006.nc wcofs_20220406_t03z_f009.nc wcofs_20220406_t03z_f012.nc wcofs_20220406_t03z_f015.nc wcofs_20220406_t03z_f018.nc wcofs_20220406_t03z_f021.nc wcofs_20220406_t03z_f024.nc wcofs_20220406_t03z_f027.nc wcofs_20220406_t03z_f030.nc wcofs_20220406_t03z_f033.nc wcofs_20220406_t03z_f036.nc wcofs_20220406_t03z_f039.nc wcofs_20220406_t03z_f042.nc wcofs_20220406_t03z_f045.nc wcofs_20220406_t03z_f048.nc wcofs_20220406_t03z_f051.nc wcofs_20220406_t03z_f054.nc wcofs_20220406_t03z_f057.nc wcofs_20220406_t03z_f060.nc wcofs_20220406_t03z_f063.nc wcofs_20220406_t03z_f066.nc wcofs_20220406_t03z_f069.nc wcofs_20220406_t03z_f072.nc" ;
}
